//
// Copyright (c) 2022 Imperas Software Ltd., www.imperas.com
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//   http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied.
//
// See the License for the specific language governing permissions and
// limitations under the License.
//
//
  
// SystemVerilog Functional Coverage Available for extensions: 
//   RV32ZCA
//   RV32ZCB
//   RV32ZCBZBB
//   RV32ZCBZMUL
//   RV32ZCMP
//   RV32ZCMT

// Uncomment to enable
//`define COVER_RV32ZCA
//`define COVER_RV32ZCB
//`define COVER_RV32ZCBZBB
//`define COVER_RV32ZCBZMUL
//`define COVER_RV32ZCMP
//`define COVER_RV32ZCMT
 

