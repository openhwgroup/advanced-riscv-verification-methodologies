//
// Copyright (c) 2022 Imperas Software Ltd., www.imperas.com
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//   http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied.
//
// See the License for the specific language governing permissions and
// limitations under the License.
//
//
 


    c_flw_cg = new(); c_flw_cg.set_inst_name("obj_c_flw");
    c_flwsp_cg = new(); c_flwsp_cg.set_inst_name("obj_c_flwsp");
    c_fsw_cg = new(); c_fsw_cg.set_inst_name("obj_c_fsw");
    c_fswsp_cg = new(); c_fswsp_cg.set_inst_name("obj_c_fswsp");


