//
// Copyright (c) 2022 Imperas Software Ltd., www.imperas.com
// 
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.0
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//   http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied.
//
// See the License for the specific language governing permissions and
// limitations under the License.
//
//
 


    fadd_s_cg = new(); fadd_s_cg.set_inst_name("obj_fadd_s");
    fclass_s_cg = new(); fclass_s_cg.set_inst_name("obj_fclass_s");
    fcvt_s_w_cg = new(); fcvt_s_w_cg.set_inst_name("obj_fcvt_s_w");
    fcvt_s_wu_cg = new(); fcvt_s_wu_cg.set_inst_name("obj_fcvt_s_wu");
    fcvt_w_s_cg = new(); fcvt_w_s_cg.set_inst_name("obj_fcvt_w_s");
    fcvt_wu_s_cg = new(); fcvt_wu_s_cg.set_inst_name("obj_fcvt_wu_s");
    fdiv_s_cg = new(); fdiv_s_cg.set_inst_name("obj_fdiv_s");
    feq_s_cg = new(); feq_s_cg.set_inst_name("obj_feq_s");
    fle_s_cg = new(); fle_s_cg.set_inst_name("obj_fle_s");
    flt_s_cg = new(); flt_s_cg.set_inst_name("obj_flt_s");
    flw_cg = new(); flw_cg.set_inst_name("obj_flw");
    fmadd_s_cg = new(); fmadd_s_cg.set_inst_name("obj_fmadd_s");
    fmax_s_cg = new(); fmax_s_cg.set_inst_name("obj_fmax_s");
    fmin_s_cg = new(); fmin_s_cg.set_inst_name("obj_fmin_s");
    fmsub_s_cg = new(); fmsub_s_cg.set_inst_name("obj_fmsub_s");
    fmul_s_cg = new(); fmul_s_cg.set_inst_name("obj_fmul_s");
    fnmadd_s_cg = new(); fnmadd_s_cg.set_inst_name("obj_fnmadd_s");
    fnmsub_s_cg = new(); fnmsub_s_cg.set_inst_name("obj_fnmsub_s");
    fsgnj_s_cg = new(); fsgnj_s_cg.set_inst_name("obj_fsgnj_s");
    fsgnjn_s_cg = new(); fsgnjn_s_cg.set_inst_name("obj_fsgnjn_s");
    fsgnjx_s_cg = new(); fsgnjx_s_cg.set_inst_name("obj_fsgnjx_s");
    fsqrt_s_cg = new(); fsqrt_s_cg.set_inst_name("obj_fsqrt_s");
    fsub_s_cg = new(); fsub_s_cg.set_inst_name("obj_fsub_s");
    fsw_cg = new(); fsw_cg.set_inst_name("obj_fsw");
    fmv_x_s_cg = new(); fmv_x_s_cg.set_inst_name("obj_fmv_x_s");
    fmv_s_x_cg = new(); fmv_s_x_cg.set_inst_name("obj_fmv_s_x");


