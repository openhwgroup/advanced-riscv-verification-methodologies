//
// Copyright (c) 2022 Imperas Software Ltd., www.imperas.com
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//   http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied.
//
// See the License for the specific language governing permissions and
// limitations under the License.
//
//
 


    cm_push_cg = new(); cm_push_cg.set_inst_name("obj_cm_push");
    cm_pop_cg = new(); cm_pop_cg.set_inst_name("obj_cm_pop");
    cm_popretz_cg = new(); cm_popretz_cg.set_inst_name("obj_cm_popretz");
    cm_popret_cg = new(); cm_popret_cg.set_inst_name("obj_cm_popret");
    cm_mvsa01_cg = new(); cm_mvsa01_cg.set_inst_name("obj_cm_mvsa01");
    cm_mva01s_cg = new(); cm_mva01s_cg.set_inst_name("obj_cm_mva01s");


