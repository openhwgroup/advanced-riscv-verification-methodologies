//
// Copyright (c) 2022 Imperas Software Ltd., www.imperas.com
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//   http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied.
//
// See the License for the specific language governing permissions and
// limitations under the License.
//
//
 


    c_add_cg = new(); c_add_cg.set_inst_name("obj_c_add");
    c_mv_cg = new(); c_mv_cg.set_inst_name("obj_c_mv");
    c_addi_cg = new(); c_addi_cg.set_inst_name("obj_c_addi");
    c_addi16sp_cg = new(); c_addi16sp_cg.set_inst_name("obj_c_addi16sp");
    c_addi4spn_cg = new(); c_addi4spn_cg.set_inst_name("obj_c_addi4spn");
    c_li_cg = new(); c_li_cg.set_inst_name("obj_c_li");
    c_lui_cg = new(); c_lui_cg.set_inst_name("obj_c_lui");
    c_and_cg = new(); c_and_cg.set_inst_name("obj_c_and");
    c_or_cg = new(); c_or_cg.set_inst_name("obj_c_or");
    c_sub_cg = new(); c_sub_cg.set_inst_name("obj_c_sub");
    c_xor_cg = new(); c_xor_cg.set_inst_name("obj_c_xor");
    c_andi_cg = new(); c_andi_cg.set_inst_name("obj_c_andi");
    c_beqz_cg = new(); c_beqz_cg.set_inst_name("obj_c_beqz");
    c_bnez_cg = new(); c_bnez_cg.set_inst_name("obj_c_bnez");
    c_j_cg = new(); c_j_cg.set_inst_name("obj_c_j");
    c_jal_cg = new(); c_jal_cg.set_inst_name("obj_c_jal");
    c_jalr_cg = new(); c_jalr_cg.set_inst_name("obj_c_jalr");
    c_jr_cg = new(); c_jr_cg.set_inst_name("obj_c_jr");
    c_lw_cg = new(); c_lw_cg.set_inst_name("obj_c_lw");
    c_lwsp_cg = new(); c_lwsp_cg.set_inst_name("obj_c_lwsp");
    c_slli_cg = new(); c_slli_cg.set_inst_name("obj_c_slli");
    c_srai_cg = new(); c_srai_cg.set_inst_name("obj_c_srai");
    c_srli_cg = new(); c_srli_cg.set_inst_name("obj_c_srli");
    c_sw_cg = new(); c_sw_cg.set_inst_name("obj_c_sw");
    c_swsp_cg = new(); c_swsp_cg.set_inst_name("obj_c_swsp");


