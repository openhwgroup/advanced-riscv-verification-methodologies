//
// Copyright (c) 2022 Imperas Software Ltd., www.imperas.com
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//   http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied.
//
// See the License for the specific language governing permissions and
// limitations under the License.
//
//
 


    c_lbu_cg = new(); c_lbu_cg.set_inst_name("obj_c_lbu");
    c_lhu_cg = new(); c_lhu_cg.set_inst_name("obj_c_lhu");
    c_lh_cg = new(); c_lh_cg.set_inst_name("obj_c_lh");
    c_sb_cg = new(); c_sb_cg.set_inst_name("obj_c_sb");
    c_sh_cg = new(); c_sh_cg.set_inst_name("obj_c_sh");
    c_zext_b_cg = new(); c_zext_b_cg.set_inst_name("obj_c_zext_b");
    c_not_cg = new(); c_not_cg.set_inst_name("obj_c_not");


