//
// Copyright (c) 2022 Imperas Software Ltd., www.imperas.com
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//   http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,
// either express or implied.
//
// See the License for the specific language governing permissions and
// limitations under the License.
//
//
 


typedef enum {
    dyn,
    rdn,
    rmm,
    rne,
    rtz,
    rup
} frm_name_t;

function frm_name_t get_frm(string s); 
    case (s)
        "rdn": return rdn;
        "rmm": return rmm;
        "rne": return rne;
        "rtz": return rtz;
        "rup": return rup;
        default: return dyn;
    endcase
endfunction


typedef struct {
    string ins_str;
    ops_t ops[6];
    int hart;
    int issue;
    bit trap;
} ins_rv32zfinx_t;


covergroup fadd_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fadd.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[3].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_frm : cross cp_fd,cp_frm  iff (ins.trap == 0) {
        option.comment = "FD FRM (ins rounding mode) Cross";
    }
    cr_fs1_frm : cross cp_fs1,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS1 FRM (ins rounding mode) Cross";
    }
    cr_fs2_frm : cross cp_fs2,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS2 FRM (ins rounding mode) Cross";
    }
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
`endif

endgroup

covergroup fclass_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fclass.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b1000000000000000000000000000000};
        bins max  = {32'b0111111111111111111111111111111};
        bins ones  = {32'b1111111111111111111111111111111};
    }
    cr_rd_fs1 : cross cp_rd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "RD FS1 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
`endif

endgroup

covergroup fcvt_s_w_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fcvt.s.w"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[2].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rs1_toggle : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_maxvals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b1000000000000000000000000000000};
        bins max  = {32'b0111111111111111111111111111111};
        bins ones  = {32'b1111111111111111111111111111111};
    }
    cr_fd_frm : cross cp_fd,cp_frm  iff (ins.trap == 0) {
        option.comment = "FD FRM (ins rounding mode) Cross";
    }
    cr_fd_rs1 : cross cp_fd,cp_rs1  iff (ins.trap == 0) {
        option.comment = "FD RS1 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
`endif

endgroup

covergroup fcvt_s_wu_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fcvt.s.wu"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_rs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "RS1 (GPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[2].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rs1_toggle : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "RS1 Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rs1_maxvals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b1000000000000000000000000000000};
        bins max  = {32'b0111111111111111111111111111111};
        bins ones  = {32'b1111111111111111111111111111111};
    }
    cr_fd_frm : cross cp_fd,cp_frm  iff (ins.trap == 0) {
        option.comment = "FD FRM (ins rounding mode) Cross";
    }
    cr_fd_rs1 : cross cp_fd,cp_rs1  iff (ins.trap == 0) {
        option.comment = "FD RS1 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
`endif

endgroup

covergroup fcvt_w_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fcvt.w.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[2].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b1000000000000000000000000000000};
        bins max  = {32'b0111111111111111111111111111111};
        bins ones  = {32'b1111111111111111111111111111111};
    }
    cr_fs1_frm : cross cp_fs1,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS1 FRM (ins rounding mode) Cross";
    }
    cr_rd_fs1 : cross cp_rd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "RD FS1 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
`endif

endgroup

covergroup fcvt_wu_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fcvt.wu.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[2].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b1000000000000000000000000000000};
        bins max  = {32'b0111111111111111111111111111111};
        bins ones  = {32'b1111111111111111111111111111111};
    }
    cr_fs1_frm : cross cp_fs1,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS1 FRM (ins rounding mode) Cross";
    }
    cr_rd_fs1 : cross cp_rd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "RD FS1 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
`endif

endgroup

covergroup fdiv_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fdiv.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[3].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_frm : cross cp_fd,cp_frm  iff (ins.trap == 0) {
        option.comment = "FD FRM (ins rounding mode) Cross";
    }
    cr_fs1_frm : cross cp_fs1,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS1 FRM (ins rounding mode) Cross";
    }
    cr_fs2_frm : cross cp_fs2,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS2 FRM (ins rounding mode) Cross";
    }
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
`endif

endgroup

covergroup feq_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "feq.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b1000000000000000000000000000000};
        bins max  = {32'b0111111111111111111111111111111};
        bins ones  = {32'b1111111111111111111111111111111};
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
    cr_rd_fs1 : cross cp_rd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "RD FS1 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
`endif

endgroup

covergroup fle_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fle.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b1000000000000000000000000000000};
        bins max  = {32'b0111111111111111111111111111111};
        bins ones  = {32'b1111111111111111111111111111111};
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
    cr_rd_fs1 : cross cp_rd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "RD FS1 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
`endif

endgroup

covergroup flt_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "flt.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_rd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "RD (GPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cp_rd_toggle : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "RD Toggle bits";
        wildcard bins bit_0_0  = {32'b???????????????????????????????0};
        wildcard bins bit_1_0  = {32'b??????????????????????????????0?};
        wildcard bins bit_2_0  = {32'b?????????????????????????????0??};
        wildcard bins bit_3_0  = {32'b????????????????????????????0???};
        wildcard bins bit_4_0  = {32'b???????????????????????????0????};
        wildcard bins bit_5_0  = {32'b??????????????????????????0?????};
        wildcard bins bit_6_0  = {32'b?????????????????????????0??????};
        wildcard bins bit_7_0  = {32'b????????????????????????0???????};
        wildcard bins bit_8_0  = {32'b???????????????????????0????????};
        wildcard bins bit_9_0  = {32'b??????????????????????0?????????};
        wildcard bins bit_10_0  = {32'b?????????????????????0??????????};
        wildcard bins bit_11_0  = {32'b????????????????????0???????????};
        wildcard bins bit_12_0  = {32'b???????????????????0????????????};
        wildcard bins bit_13_0  = {32'b??????????????????0?????????????};
        wildcard bins bit_14_0  = {32'b?????????????????0??????????????};
        wildcard bins bit_15_0  = {32'b????????????????0???????????????};
        wildcard bins bit_16_0  = {32'b???????????????0????????????????};
        wildcard bins bit_17_0  = {32'b??????????????0?????????????????};
        wildcard bins bit_18_0  = {32'b?????????????0??????????????????};
        wildcard bins bit_19_0  = {32'b????????????0???????????????????};
        wildcard bins bit_20_0  = {32'b???????????0????????????????????};
        wildcard bins bit_21_0  = {32'b??????????0?????????????????????};
        wildcard bins bit_22_0  = {32'b?????????0??????????????????????};
        wildcard bins bit_23_0  = {32'b????????0???????????????????????};
        wildcard bins bit_24_0  = {32'b???????0????????????????????????};
        wildcard bins bit_25_0  = {32'b??????0?????????????????????????};
        wildcard bins bit_26_0  = {32'b?????0??????????????????????????};
        wildcard bins bit_27_0  = {32'b????0???????????????????????????};
        wildcard bins bit_28_0  = {32'b???0????????????????????????????};
        wildcard bins bit_29_0  = {32'b??0?????????????????????????????};
        wildcard bins bit_30_0  = {32'b?0??????????????????????????????};
        wildcard bins bit_31_0  = {32'b0???????????????????????????????};
        wildcard bins bit_0_1  = {32'b???????????????????????????????1};
        wildcard bins bit_1_1  = {32'b??????????????????????????????1?};
        wildcard bins bit_2_1  = {32'b?????????????????????????????1??};
        wildcard bins bit_3_1  = {32'b????????????????????????????1???};
        wildcard bins bit_4_1  = {32'b???????????????????????????1????};
        wildcard bins bit_5_1  = {32'b??????????????????????????1?????};
        wildcard bins bit_6_1  = {32'b?????????????????????????1??????};
        wildcard bins bit_7_1  = {32'b????????????????????????1???????};
        wildcard bins bit_8_1  = {32'b???????????????????????1????????};
        wildcard bins bit_9_1  = {32'b??????????????????????1?????????};
        wildcard bins bit_10_1  = {32'b?????????????????????1??????????};
        wildcard bins bit_11_1  = {32'b????????????????????1???????????};
        wildcard bins bit_12_1  = {32'b???????????????????1????????????};
        wildcard bins bit_13_1  = {32'b??????????????????1?????????????};
        wildcard bins bit_14_1  = {32'b?????????????????1??????????????};
        wildcard bins bit_15_1  = {32'b????????????????1???????????????};
        wildcard bins bit_16_1  = {32'b???????????????1????????????????};
        wildcard bins bit_17_1  = {32'b??????????????1?????????????????};
        wildcard bins bit_18_1  = {32'b?????????????1??????????????????};
        wildcard bins bit_19_1  = {32'b????????????1???????????????????};
        wildcard bins bit_20_1  = {32'b???????????1????????????????????};
        wildcard bins bit_21_1  = {32'b??????????1?????????????????????};
        wildcard bins bit_22_1  = {32'b?????????1??????????????????????};
        wildcard bins bit_23_1  = {32'b????????1???????????????????????};
        wildcard bins bit_24_1  = {32'b???????1????????????????????????};
        wildcard bins bit_25_1  = {32'b??????1?????????????????????????};
        wildcard bins bit_26_1  = {32'b?????1??????????????????????????};
        wildcard bins bit_27_1  = {32'b????1???????????????????????????};
        wildcard bins bit_28_1  = {32'b???1????????????????????????????};
        wildcard bins bit_29_1  = {32'b??1?????????????????????????????};
        wildcard bins bit_30_1  = {32'b?1??????????????????????????????};
        wildcard bins bit_31_1  = {32'b1???????????????????????????????};
    }
    cp_rd_maxvals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "RD Max values";
        bins zeros  = {0};
        bins min  = {32'b1000000000000000000000000000000};
        bins max  = {32'b0111111111111111111111111111111};
        bins ones  = {32'b1111111111111111111111111111111};
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
    cr_rd_fs1 : cross cp_rd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "RD FS1 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
`endif

endgroup

covergroup fmadd_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fmadd.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }
    cp_fs3 : coverpoint get_gpr_reg(ins.ops[3].key)  iff (ins.trap == 0) {
        option.comment = "FS3 (FPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[4].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_frm : cross cp_fd,cp_frm  iff (ins.trap == 0) {
        option.comment = "FD FRM (ins rounding mode) Cross";
    }
    cr_fs1_frm : cross cp_fs1,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS1 FRM (ins rounding mode) Cross";
    }
    cr_fs2_frm : cross cp_fs2,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS2 FRM (ins rounding mode) Cross";
    }
    cr_fs3_frm : cross cp_fs3,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS3 FRM (ins rounding mode) Cross";
    }
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fd_fs3 : cross cp_fd,cp_fs3  iff (ins.trap == 0) {
        option.comment = "FD FS3 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
    cr_fs1_fs2_fs3 : cross cp_fs1,cp_fs2,cp_fs3  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 FS3 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs3_vals : coverpoint unsigned'(int'(ins.ops[3].val))  iff (ins.trap == 0) {
        option.comment = "FS3 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
    cr_fs3_vals : cross cp_fs3,cp_fs3_vals  iff (ins.trap == 0) {
        option.comment = "FS3 FPU values Cross";
    }
`endif

endgroup

covergroup fmax_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fmax.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
`endif

endgroup

covergroup fmin_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fmin.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
`endif

endgroup

covergroup fmsub_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fmsub.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }
    cp_fs3 : coverpoint get_gpr_reg(ins.ops[3].key)  iff (ins.trap == 0) {
        option.comment = "FS3 (FPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[4].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_frm : cross cp_fd,cp_frm  iff (ins.trap == 0) {
        option.comment = "FD FRM (ins rounding mode) Cross";
    }
    cr_fs1_frm : cross cp_fs1,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS1 FRM (ins rounding mode) Cross";
    }
    cr_fs2_frm : cross cp_fs2,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS2 FRM (ins rounding mode) Cross";
    }
    cr_fs3_frm : cross cp_fs3,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS3 FRM (ins rounding mode) Cross";
    }
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fd_fs3 : cross cp_fd,cp_fs3  iff (ins.trap == 0) {
        option.comment = "FD FS3 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
    cr_fs1_fs2_fs3 : cross cp_fs1,cp_fs2,cp_fs3  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 FS3 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs3_vals : coverpoint unsigned'(int'(ins.ops[3].val))  iff (ins.trap == 0) {
        option.comment = "FS3 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
    cr_fs3_vals : cross cp_fs3,cp_fs3_vals  iff (ins.trap == 0) {
        option.comment = "FS3 FPU values Cross";
    }
`endif

endgroup

covergroup fmul_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fmul.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[3].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_frm : cross cp_fd,cp_frm  iff (ins.trap == 0) {
        option.comment = "FD FRM (ins rounding mode) Cross";
    }
    cr_fs1_frm : cross cp_fs1,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS1 FRM (ins rounding mode) Cross";
    }
    cr_fs2_frm : cross cp_fs2,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS2 FRM (ins rounding mode) Cross";
    }
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
`endif

endgroup

covergroup fnmadd_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fnmadd.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }
    cp_fs3 : coverpoint get_gpr_reg(ins.ops[3].key)  iff (ins.trap == 0) {
        option.comment = "FS3 (FPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[4].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_frm : cross cp_fd,cp_frm  iff (ins.trap == 0) {
        option.comment = "FD FRM (ins rounding mode) Cross";
    }
    cr_fs1_frm : cross cp_fs1,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS1 FRM (ins rounding mode) Cross";
    }
    cr_fs2_frm : cross cp_fs2,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS2 FRM (ins rounding mode) Cross";
    }
    cr_fs3_frm : cross cp_fs3,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS3 FRM (ins rounding mode) Cross";
    }
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fd_fs3 : cross cp_fd,cp_fs3  iff (ins.trap == 0) {
        option.comment = "FD FS3 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
    cr_fs1_fs2_fs3 : cross cp_fs1,cp_fs2,cp_fs3  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 FS3 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs3_vals : coverpoint unsigned'(int'(ins.ops[3].val))  iff (ins.trap == 0) {
        option.comment = "FS3 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
    cr_fs3_vals : cross cp_fs3,cp_fs3_vals  iff (ins.trap == 0) {
        option.comment = "FS3 FPU values Cross";
    }
`endif

endgroup

covergroup fnmsub_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fnmsub.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }
    cp_fs3 : coverpoint get_gpr_reg(ins.ops[3].key)  iff (ins.trap == 0) {
        option.comment = "FS3 (FPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[4].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_frm : cross cp_fd,cp_frm  iff (ins.trap == 0) {
        option.comment = "FD FRM (ins rounding mode) Cross";
    }
    cr_fs1_frm : cross cp_fs1,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS1 FRM (ins rounding mode) Cross";
    }
    cr_fs2_frm : cross cp_fs2,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS2 FRM (ins rounding mode) Cross";
    }
    cr_fs3_frm : cross cp_fs3,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS3 FRM (ins rounding mode) Cross";
    }
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fd_fs3 : cross cp_fd,cp_fs3  iff (ins.trap == 0) {
        option.comment = "FD FS3 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
    cr_fs1_fs2_fs3 : cross cp_fs1,cp_fs2,cp_fs3  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 FS3 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs3_vals : coverpoint unsigned'(int'(ins.ops[3].val))  iff (ins.trap == 0) {
        option.comment = "FS3 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
    cr_fs3_vals : cross cp_fs3,cp_fs3_vals  iff (ins.trap == 0) {
        option.comment = "FS3 FPU values Cross";
    }
`endif

endgroup

covergroup fsgnj_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fsgnj.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
`endif

endgroup

covergroup fsgnjn_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fsgnjn.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
`endif

endgroup

covergroup fsgnjx_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fsgnjx.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
`endif

endgroup

covergroup fsqrt_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fsqrt.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[2].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_frm : cross cp_fd,cp_frm  iff (ins.trap == 0) {
        option.comment = "FD FRM (ins rounding mode) Cross";
    }
    cr_fs1_frm : cross cp_fs1,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS1 FRM (ins rounding mode) Cross";
    }
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
`endif

endgroup

covergroup fsub_s_cg with function sample(ins_rv32zfinx_t ins);
    option.per_instance = 1; 
    cp_asm_count : coverpoint ins.ins_str == "fsub.s"  iff (ins.trap == 0) {
        option.comment = "Number of times instruction is executed";
        bins count[]  = {1};
    }
    cp_fd : coverpoint get_gpr_reg(ins.ops[0].key)  iff (ins.trap == 0) {
        option.comment = "FD (FPR) register assignment";
    }
    cp_fs1 : coverpoint get_gpr_reg(ins.ops[1].key)  iff (ins.trap == 0) {
        option.comment = "FS1 (FPR) register assignment";
    }
    cp_fs2 : coverpoint get_gpr_reg(ins.ops[2].key)  iff (ins.trap == 0) {
        option.comment = "FS2 (FPR) register assignment";
    }
    cp_frm : coverpoint get_frm(ins.ops[3].val)  iff (ins.trap == 0) {
        option.comment = "Floating Point FRM (Rounding mode) given as an operand";
    }
    cp_csr_fcsr_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "fcsr", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fcsr_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fcsr", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fcsr CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }
    cp_csr_frm_frm : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_BEFORE, "frm", "frm")  iff (ins.trap == 0) {
        option.comment = "Value of frm CSR, frm field";
        bins rne  = {3'b000};
        bins rtz  = {3'b001};
        bins rdn  = {3'b010};
        bins rup  = {3'b011};
        bins rmm  = {3'b100};
        bins illegal  = default;
    }
    cp_csr_fflags_fflags : coverpoint get_csr_val(ins.hart, ins.issue, `SAMPLE_AFTER, "fflags", "fflags")  iff (ins.trap == 0) {
        option.comment = "Value of fflags CSR, fflags field";
        wildcard bins NX  = {5'b????1};
        wildcard bins UF  = {5'b???1?};
        wildcard bins OF  = {5'b??1??};
        wildcard bins DZ  = {5'b?1???};
        wildcard bins NV  = {5'b1????};
    }

`ifdef COVER_LEVEL_COMPL_EXT
    cr_fd_frm : cross cp_fd,cp_frm  iff (ins.trap == 0) {
        option.comment = "FD FRM (ins rounding mode) Cross";
    }
    cr_fs1_frm : cross cp_fs1,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS1 FRM (ins rounding mode) Cross";
    }
    cr_fs2_frm : cross cp_fs2,cp_frm  iff (ins.trap == 0) {
        option.comment = "FS2 FRM (ins rounding mode) Cross";
    }
    cr_fd_fs1 : cross cp_fd,cp_fs1  iff (ins.trap == 0) {
        option.comment = "FD FS1 Cross";
    }
    cr_fd_fs2 : cross cp_fd,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FD FS2 Cross";
    }
    cr_fs1_fs2 : cross cp_fs1,cp_fs2  iff (ins.trap == 0) {
        option.comment = "FS1 FS2 Cross";
    }
`endif


`ifdef COVER_LEVEL_DV_UP_BAS
    cp_fd_vals : coverpoint unsigned'(int'(ins.ops[0].val))  iff (ins.trap == 0) {
        option.comment = "FD FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs1_vals : coverpoint unsigned'(int'(ins.ops[1].val))  iff (ins.trap == 0) {
        option.comment = "FS1 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cp_fs2_vals : coverpoint unsigned'(int'(ins.ops[2].val))  iff (ins.trap == 0) {
        option.comment = "FS2 FPU Special values";
        bins plus_0p0  = {32'h0};
        bins minus_0p0  = {32'h80000000};
        bins plus_minnorm  = {32'h800000};
        bins minus_minnorm  = {32'h80800000};
        bins plus_minnorm_div2  = {32'h400000};
        bins minus_minnorm_div2  = {32'h80400000};
        bins plus_maxnorm  = {32'h7f7fffff};
        bins minus_maxnorm  = {32'hff7fffff};
        bins plus_max_subnorm  = {32'h7fffff};
        bins minus_max_subnorm  = {32'h807fffff};
        bins plus_min_subnorm  = {32'h1};
        bins minus_min_subnorm  = {32'h80000001};
        bins plus_infinity  = {32'h7f800000};
        bins minus_infinity  = {32'hff800000};
        bins plus_QNaN  = {32'h7fc12345};
    }
    cr_fd_vals : cross cp_fd,cp_fd_vals  iff (ins.trap == 0) {
        option.comment = "FD FPU values Cross";
    }
    cr_fs1_vals : cross cp_fs1,cp_fs1_vals  iff (ins.trap == 0) {
        option.comment = "FS1 FPU values Cross";
    }
    cr_fs2_vals : cross cp_fs2,cp_fs2_vals  iff (ins.trap == 0) {
        option.comment = "FS2 FPU values Cross";
    }
`endif

endgroup


function ins_rv32zfinx_t get_rv32zfinx_inst(bit trap, int hart, int issue, string disass); // break and move this first bit out
    string insbin, ins_str, op[6], key, val;
    ins_rv32zfinx_t ins;
    int num, i, j;
    string s = disass;
    foreach (disass[c]) begin
        s[c] = (disass[c] == ",")? " " : disass[c];
    end
    ins.hart = hart;
    ins.issue = issue;
    ins.trap = trap;
    num = $sscanf (s, "%s %s %s %s %s %s %s %s", insbin, ins_str, op[0], op[1], op[2], op[3], op[4], op[5]);
    ins.ins_str = ins_str;
    for (i=0; i<num-2; i++) begin
        key = op[i];
        ins.ops[i].key=op[i]; // in case we dont update it as an indexed
        ins.ops[i].val=""; // not used
        for (j = 0; j < key.len(); j++) begin // if indexed addressing, convert offset(rs1) to op[i].key=rs1 op[i+1].key=offset
            if (key[j] == "(") begin
                ins.ops[i].key = key.substr(0,j-1); // offset
                ins.ops[i+1].key = key.substr(j+1,key.len()-2);
                i++; // step over +1
                //$display("indirect ins_str(%s) op[0](%0s).key(%s) op[1](%s).key(%s) op[2](%s).key(%s) op[3](%s).key(%s)", 
                //    ins_str, op[0], ins.ops[0].key, op[1], ins.ops[1].key, op[2], ins.ops[2].key, op[3], ins.ops[3].key);
                break;
            end
        end
    end
    for (i=0; i<num-2; i++) begin
        if (ins.ops[i].key[0] == "x") begin
            int idx = get_gpr_num(ins.ops[i].key);
            //$display("SAMPLE: %0s op[%0d]=%0s gpr(%0d)", ins_str,i, ins.ops[i].key, idx);
            if (idx < 0) begin
                ins.ops[i].val = ins.ops[i].key; // it is an immed already there
            end else begin
                ins.ops[i].val = string'(this.rvvi.x_wdata[hart][issue][idx]);
            end
        end else if (ins.ops[i].key[0] == "f") begin
            int idx = get_fpr_num(ins.ops[i].key);
            if (idx < 0) begin
                ins.ops[i].val = ins.ops[i].key; // it is an immed already there
            end else begin
                ins.ops[i].val = string'(this.rvvi.f_wdata[hart][issue][idx]);
            end
        end else begin
            ins.ops[i].val = ins.ops[i].key;
        end       
    end
    return ins;
endfunction

function void rv32zfinx_sample(string inst_name, bit trap, int hart, int issue, string disass);
    case (inst_name)
        "fadd.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fadd_s_cg.sample(ins); end
        "fclass.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fclass_s_cg.sample(ins); end
        "fcvt.s.w"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fcvt_s_w_cg.sample(ins); end
        "fcvt.s.wu"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fcvt_s_wu_cg.sample(ins); end
        "fcvt.w.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fcvt_w_s_cg.sample(ins); end
        "fcvt.wu.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fcvt_wu_s_cg.sample(ins); end
        "fdiv.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fdiv_s_cg.sample(ins); end
        "feq.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); feq_s_cg.sample(ins); end
        "fle.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fle_s_cg.sample(ins); end
        "flt.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); flt_s_cg.sample(ins); end
        "fmadd.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fmadd_s_cg.sample(ins); end
        "fmax.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fmax_s_cg.sample(ins); end
        "fmin.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fmin_s_cg.sample(ins); end
        "fmsub.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fmsub_s_cg.sample(ins); end
        "fmul.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fmul_s_cg.sample(ins); end
        "fnmadd.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fnmadd_s_cg.sample(ins); end
        "fnmsub.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fnmsub_s_cg.sample(ins); end
        "fsgnj.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fsgnj_s_cg.sample(ins); end
        "fsgnjn.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fsgnjn_s_cg.sample(ins); end
        "fsgnjx.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fsgnjx_s_cg.sample(ins); end
        "fsqrt.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fsqrt_s_cg.sample(ins); end
        "fsub.s"     : begin ins_rv32zfinx_t ins = get_rv32zfinx_inst(trap, hart, issue, disass); fsub_s_cg.sample(ins); end
    endcase
endfunction


